//ld_op.v, 32-bit LOAD DIRECT instruction module 

`timescale 1ns/10ps

module ld_op (
);
