//mfhi_op.v, 32-bit MOVE FROM HI instruction module 

`timescale 1ns/10ps

module mfhi_op (
);
