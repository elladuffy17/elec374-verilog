/* also for the bus we need a 32-to-5 encoder, which is a combinational circuit. 
It has 2^n input lines and n output lines. It takes up these 2^n input data and encodes them into n-bit data. 
Therefore, it produces the binary code equivalent of the input line, which is active high */

module encoder(
  output reg [4:0] output,
  input [31:0] input);

  always @(input)
  begin
    case (input)
      'b00000000000000000000000000000001 : out <= 'b00000; //32 bit input to a 4 bit output
      'b00000000000000000000000000000010 : out <= 'b00001;
      'b00000000000000000000000000000100 : out <= 'b00010;
      'b00000000000000000000000000001000 : out <= 'b00011;
      'b00000000000000000000000000010000 : out <= 'b00100;
      'b00000000000000000000000000100000 : out <= 'b00101;
      'b00000000000000000000000001000000 : out <= 'b00110;
      'b00000000000000000000000010000000 : out <= 'b00111;
      'b00000000000000000000000100000000 : out <= 'b01000;
      'b00000000000000000000001000000000 : out <= 'b01001;
      'b00000000000000000000010000000000 : out <= 'b01010;
      'b00000000000000000000100000000000 : out <= 'b01011;
      'b00000000000000000001000000000000 : out <= 'b01100;
      'b00000000000000000010000000000000 : out <= 'b01101;
      'b00000000000000000100000000000000 : out <= 'b01110;
      'b00000000000000001000000000000000 : out <= 'b01111;
      'b00000000000000010000000000000000 : out <= 'b10000;
      'b00000000000000100000000000000000 : out <= 'b10001;
      'b00000000000001000000000000000000 : out <= 'b10010;
      'b00000000000010000000000000000000 : out <= 'b10011;
      'b00000000000100000000000000000000 : out <= 'b10100;
      'b00000000001000000000000000000000 : out <= 'b10101;
      'b00000000010000000000000000000000 : out <= 'b10110;
      'b00000000100000000000000000000000 : out <= 'b10111;
      'b00000001000000000000000000000000 : out <= 'b11000;
      'b00000010000000000000000000000000 : out <= 'b11001;
      'b00000100000000000000000000000000 : out <= 'b11010;
      'b00001000000000000000000000000000 : out <= 'b11011;
      'b00010000000000000000000000000000 : out <= 'b11100;
      'b00100000000000000000000000000000 : out <= 'b11101;
      'b01000000000000000000000000000000 : out <= 'b11110;
      'b10000000000000000000000000000000 : out <= 'b11111;
    default: out <= 0;
      
  endcase

  end
endmodule
