//out_op.v, 32-bit OUTPUT instruction module 

`timescale 1ns/10ps

module out_op (
);
