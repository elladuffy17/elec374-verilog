//ori_op.v, 32-bit OR IMMEDIATE instruction module 

`timescale 1ns/10ps

module ori_op (
);
