//out_op.v, 32-bit OUT instruction module 

`timescale 1ns/10ps

module out_op (
);
