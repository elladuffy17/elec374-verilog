//branch_instr_tb.v, testbench for the BRANCH INSTRUCTIONS (brzr, brnz, brpl, brmi)

`timescale 1ns/10ps

module branch_instr_tb;

endmodule
