module CONFFLogic ();
