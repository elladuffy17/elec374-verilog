//andi_op.v, 32-bit AND IMMEDIATE instruction module 

`timescale 1ns/10ps

module andi_op (
);
