//mflo_op.v, 32-bit MOVE FROM LO instruction module 

`timescale 1ns/10ps

module mflo_op (
);
