//jal_op.v, 32-bit JUMP AND LINK instruction module 

`timescale 1ns/10ps

module jal_op (
);
