//ldi_op.v, 32-bit LOAD IMMEDIATE instruction module 

`timescale 1ns/10ps

module ldi_op (
);
