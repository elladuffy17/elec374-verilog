//jr_op.v, 32-bit RETURN FROM PROCEDURE instruction module 

`timescale 1ns/10ps

module jr_op (
);
