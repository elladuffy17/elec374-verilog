//st_op.v, 32-bit STORE DIRECT instruction module 

`timescale 1ns/10ps

module st_op (
);
