//in_op.v, 32-bit INPUT instruction module 

`timescale 1ns/10ps

module in_op (
);
