//addi_op.v, 32-bit ADD IMMEDIATE instruction module 

`timescale 1ns/10ps

module addi_op (
);
